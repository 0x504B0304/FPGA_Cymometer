
module issp (
	source,
	probe);	

	output	[22:0]	source;
	input	[63:0]	probe;
endmodule
